`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: VIT
// Engineer: Rohan Boge
//////////////////////////////////////////////////////////////////////////////////
module FA(a,b,cin,sum,carry);	input a,b,cin;
	output sum,carry;
	
	assign sum = a^b^cin;
	assign carry = (a&b) | (b&cin) | (a&cin);

endmodule
